library verilog;
use verilog.vl_types.all;
entity SDB_tb is
end SDB_tb;
